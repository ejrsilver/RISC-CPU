// This adder is only used for the CSA, which is why I used Add_Generator.java 
// to create the logic instead of combining modules. Honestly 
// it's just funnier but might technically be faster as well, who knows!
module add_64(
    input [63:0] A, B,
    input Cin,
    output [63:0] Z,
    output Cout);

    wire [63:0] P,G,c;
    assign P = A^B; 
    assign G = A&B;
    assign c[0] = Cin;
assign c[1] = G[0] | (P[0]&c[0]);
assign c[2] = G[1] | (P[1]&G[0]) | (P[1]&P[0]&c[0]);
assign c[3] = G[2] | (P[2]&G[1]) | (P[2]&P[1]&G[0]) | (P[2]&P[1]&P[0]&c[0]);
assign c[4] = G[3] | (P[3]&G[2]) | (P[3]&P[2]&G[1]) | (P[3]&P[2]&P[1]&G[0]) | (P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[5] = G[4] | (P[4]&G[3]) | (P[4]&P[3]&G[2]) | (P[4]&P[3]&P[2]&G[1]) | (P[4]&P[3]&P[2]&P[1]&G[0]) | (P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[6] = G[5] | (P[5]&G[4]) | (P[5]&P[4]&G[3]) | (P[5]&P[4]&P[3]&G[2]) | (P[5]&P[4]&P[3]&P[2]&G[1]) | (P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[7] = G[6] | (P[6]&G[5]) | (P[6]&P[5]&G[4]) | (P[6]&P[5]&P[4]&G[3]) | (P[6]&P[5]&P[4]&P[3]&G[2]) | (P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[8] = G[7] | (P[7]&G[6]) | (P[7]&P[6]&G[5]) | (P[7]&P[6]&P[5]&G[4]) | (P[7]&P[6]&P[5]&P[4]&G[3]) | (P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[9] = G[8] | (P[8]&G[7]) | (P[8]&P[7]&G[6]) | (P[8]&P[7]&P[6]&G[5]) | (P[8]&P[7]&P[6]&P[5]&G[4]) | (P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[10] = G[9] | (P[9]&G[8]) | (P[9]&P[8]&G[7]) | (P[9]&P[8]&P[7]&G[6]) | (P[9]&P[8]&P[7]&P[6]&G[5]) | (P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[11] = G[10] | (P[10]&G[9]) | (P[10]&P[9]&G[8]) | (P[10]&P[9]&P[8]&G[7]) | (P[10]&P[9]&P[8]&P[7]&G[6]) | (P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[12] = G[11] | (P[11]&G[10]) | (P[11]&P[10]&G[9]) | (P[11]&P[10]&P[9]&G[8]) | (P[11]&P[10]&P[9]&P[8]&G[7]) | (P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[13] = G[12] | (P[12]&G[11]) | (P[12]&P[11]&G[10]) | (P[12]&P[11]&P[10]&G[9]) | (P[12]&P[11]&P[10]&P[9]&G[8]) | (P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[14] = G[13] | (P[13]&G[12]) | (P[13]&P[12]&G[11]) | (P[13]&P[12]&P[11]&G[10]) | (P[13]&P[12]&P[11]&P[10]&G[9]) | (P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[15] = G[14] | (P[14]&G[13]) | (P[14]&P[13]&G[12]) | (P[14]&P[13]&P[12]&G[11]) | (P[14]&P[13]&P[12]&P[11]&G[10]) | (P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[16] = G[15] | (P[15]&G[14]) | (P[15]&P[14]&G[13]) | (P[15]&P[14]&P[13]&G[12]) | (P[15]&P[14]&P[13]&P[12]&G[11]) | (P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[17] = G[16] | (P[16]&G[15]) | (P[16]&P[15]&G[14]) | (P[16]&P[15]&P[14]&G[13]) | (P[16]&P[15]&P[14]&P[13]&G[12]) | (P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[18] = G[17] | (P[17]&G[16]) | (P[17]&P[16]&G[15]) | (P[17]&P[16]&P[15]&G[14]) | (P[17]&P[16]&P[15]&P[14]&G[13]) | (P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[19] = G[18] | (P[18]&G[17]) | (P[18]&P[17]&G[16]) | (P[18]&P[17]&P[16]&G[15]) | (P[18]&P[17]&P[16]&P[15]&G[14]) | (P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[20] = G[19] | (P[19]&G[18]) | (P[19]&P[18]&G[17]) | (P[19]&P[18]&P[17]&G[16]) | (P[19]&P[18]&P[17]&P[16]&G[15]) | (P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[21] = G[20] | (P[20]&G[19]) | (P[20]&P[19]&G[18]) | (P[20]&P[19]&P[18]&G[17]) | (P[20]&P[19]&P[18]&P[17]&G[16]) | (P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[22] = G[21] | (P[21]&G[20]) | (P[21]&P[20]&G[19]) | (P[21]&P[20]&P[19]&G[18]) | (P[21]&P[20]&P[19]&P[18]&G[17]) | (P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[23] = G[22] | (P[22]&G[21]) | (P[22]&P[21]&G[20]) | (P[22]&P[21]&P[20]&G[19]) | (P[22]&P[21]&P[20]&P[19]&G[18]) | (P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[24] = G[23] | (P[23]&G[22]) | (P[23]&P[22]&G[21]) | (P[23]&P[22]&P[21]&G[20]) | (P[23]&P[22]&P[21]&P[20]&G[19]) | (P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[25] = G[24] | (P[24]&G[23]) | (P[24]&P[23]&G[22]) | (P[24]&P[23]&P[22]&G[21]) | (P[24]&P[23]&P[22]&P[21]&G[20]) | (P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[26] = G[25] | (P[25]&G[24]) | (P[25]&P[24]&G[23]) | (P[25]&P[24]&P[23]&G[22]) | (P[25]&P[24]&P[23]&P[22]&G[21]) | (P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[27] = G[26] | (P[26]&G[25]) | (P[26]&P[25]&G[24]) | (P[26]&P[25]&P[24]&G[23]) | (P[26]&P[25]&P[24]&P[23]&G[22]) | (P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[28] = G[27] | (P[27]&G[26]) | (P[27]&P[26]&G[25]) | (P[27]&P[26]&P[25]&G[24]) | (P[27]&P[26]&P[25]&P[24]&G[23]) | (P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[29] = G[28] | (P[28]&G[27]) | (P[28]&P[27]&G[26]) | (P[28]&P[27]&P[26]&G[25]) | (P[28]&P[27]&P[26]&P[25]&G[24]) | (P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[30] = G[29] | (P[29]&G[28]) | (P[29]&P[28]&G[27]) | (P[29]&P[28]&P[27]&G[26]) | (P[29]&P[28]&P[27]&P[26]&G[25]) | (P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[31] = G[30] | (P[30]&G[29]) | (P[30]&P[29]&G[28]) | (P[30]&P[29]&P[28]&G[27]) | (P[30]&P[29]&P[28]&P[27]&G[26]) | (P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[32] = G[31] | (P[31]&G[30]) | (P[31]&P[30]&G[29]) | (P[31]&P[30]&P[29]&G[28]) | (P[31]&P[30]&P[29]&P[28]&G[27]) | (P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[33] = G[32] | (P[32]&G[31]) | (P[32]&P[31]&G[30]) | (P[32]&P[31]&P[30]&G[29]) | (P[32]&P[31]&P[30]&P[29]&G[28]) | (P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[34] = G[33] | (P[33]&G[32]) | (P[33]&P[32]&G[31]) | (P[33]&P[32]&P[31]&G[30]) | (P[33]&P[32]&P[31]&P[30]&G[29]) | (P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[35] = G[34] | (P[34]&G[33]) | (P[34]&P[33]&G[32]) | (P[34]&P[33]&P[32]&G[31]) | (P[34]&P[33]&P[32]&P[31]&G[30]) | (P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[36] = G[35] | (P[35]&G[34]) | (P[35]&P[34]&G[33]) | (P[35]&P[34]&P[33]&G[32]) | (P[35]&P[34]&P[33]&P[32]&G[31]) | (P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[37] = G[36] | (P[36]&G[35]) | (P[36]&P[35]&G[34]) | (P[36]&P[35]&P[34]&G[33]) | (P[36]&P[35]&P[34]&P[33]&G[32]) | (P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[38] = G[37] | (P[37]&G[36]) | (P[37]&P[36]&G[35]) | (P[37]&P[36]&P[35]&G[34]) | (P[37]&P[36]&P[35]&P[34]&G[33]) | (P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[39] = G[38] | (P[38]&G[37]) | (P[38]&P[37]&G[36]) | (P[38]&P[37]&P[36]&G[35]) | (P[38]&P[37]&P[36]&P[35]&G[34]) | (P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[40] = G[39] | (P[39]&G[38]) | (P[39]&P[38]&G[37]) | (P[39]&P[38]&P[37]&G[36]) | (P[39]&P[38]&P[37]&P[36]&G[35]) | (P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[41] = G[40] | (P[40]&G[39]) | (P[40]&P[39]&G[38]) | (P[40]&P[39]&P[38]&G[37]) | (P[40]&P[39]&P[38]&P[37]&G[36]) | (P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[42] = G[41] | (P[41]&G[40]) | (P[41]&P[40]&G[39]) | (P[41]&P[40]&P[39]&G[38]) | (P[41]&P[40]&P[39]&P[38]&G[37]) | (P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[43] = G[42] | (P[42]&G[41]) | (P[42]&P[41]&G[40]) | (P[42]&P[41]&P[40]&G[39]) | (P[42]&P[41]&P[40]&P[39]&G[38]) | (P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[44] = G[43] | (P[43]&G[42]) | (P[43]&P[42]&G[41]) | (P[43]&P[42]&P[41]&G[40]) | (P[43]&P[42]&P[41]&P[40]&G[39]) | (P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[45] = G[44] | (P[44]&G[43]) | (P[44]&P[43]&G[42]) | (P[44]&P[43]&P[42]&G[41]) | (P[44]&P[43]&P[42]&P[41]&G[40]) | (P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[46] = G[45] | (P[45]&G[44]) | (P[45]&P[44]&G[43]) | (P[45]&P[44]&P[43]&G[42]) | (P[45]&P[44]&P[43]&P[42]&G[41]) | (P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[47] = G[46] | (P[46]&G[45]) | (P[46]&P[45]&G[44]) | (P[46]&P[45]&P[44]&G[43]) | (P[46]&P[45]&P[44]&P[43]&G[42]) | (P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[48] = G[47] | (P[47]&G[46]) | (P[47]&P[46]&G[45]) | (P[47]&P[46]&P[45]&G[44]) | (P[47]&P[46]&P[45]&P[44]&G[43]) | (P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[49] = G[48] | (P[48]&G[47]) | (P[48]&P[47]&G[46]) | (P[48]&P[47]&P[46]&G[45]) | (P[48]&P[47]&P[46]&P[45]&G[44]) | (P[48]&P[47]&P[46]&P[45]&P[44]&G[43]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[50] = G[49] | (P[49]&G[48]) | (P[49]&P[48]&G[47]) | (P[49]&P[48]&P[47]&G[46]) | (P[49]&P[48]&P[47]&P[46]&G[45]) | (P[49]&P[48]&P[47]&P[46]&P[45]&G[44]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&G[43]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[51] = G[50] | (P[50]&G[49]) | (P[50]&P[49]&G[48]) | (P[50]&P[49]&P[48]&G[47]) | (P[50]&P[49]&P[48]&P[47]&G[46]) | (P[50]&P[49]&P[48]&P[47]&P[46]&G[45]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&G[44]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&G[43]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[52] = G[51] | (P[51]&G[50]) | (P[51]&P[50]&G[49]) | (P[51]&P[50]&P[49]&G[48]) | (P[51]&P[50]&P[49]&P[48]&G[47]) | (P[51]&P[50]&P[49]&P[48]&P[47]&G[46]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&G[45]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&G[44]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&G[43]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[53] = G[52] | (P[52]&G[51]) | (P[52]&P[51]&G[50]) | (P[52]&P[51]&P[50]&G[49]) | (P[52]&P[51]&P[50]&P[49]&G[48]) | (P[52]&P[51]&P[50]&P[49]&P[48]&G[47]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&G[46]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&G[45]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&G[44]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&G[43]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[54] = G[53] | (P[53]&G[52]) | (P[53]&P[52]&G[51]) | (P[53]&P[52]&P[51]&G[50]) | (P[53]&P[52]&P[51]&P[50]&G[49]) | (P[53]&P[52]&P[51]&P[50]&P[49]&G[48]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&G[47]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&G[46]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&G[45]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&G[44]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&G[43]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[55] = G[54] | (P[54]&G[53]) | (P[54]&P[53]&G[52]) | (P[54]&P[53]&P[52]&G[51]) | (P[54]&P[53]&P[52]&P[51]&G[50]) | (P[54]&P[53]&P[52]&P[51]&P[50]&G[49]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&G[48]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&G[47]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&G[46]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&G[45]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&G[44]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&G[43]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[56] = G[55] | (P[55]&G[54]) | (P[55]&P[54]&G[53]) | (P[55]&P[54]&P[53]&G[52]) | (P[55]&P[54]&P[53]&P[52]&G[51]) | (P[55]&P[54]&P[53]&P[52]&P[51]&G[50]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&G[49]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&G[48]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&G[47]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&G[46]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&G[45]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&G[44]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&G[43]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[57] = G[56] | (P[56]&G[55]) | (P[56]&P[55]&G[54]) | (P[56]&P[55]&P[54]&G[53]) | (P[56]&P[55]&P[54]&P[53]&G[52]) | (P[56]&P[55]&P[54]&P[53]&P[52]&G[51]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&G[50]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&G[49]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&G[48]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&G[47]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&G[46]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&G[45]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&G[44]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&G[43]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[58] = G[57] | (P[57]&G[56]) | (P[57]&P[56]&G[55]) | (P[57]&P[56]&P[55]&G[54]) | (P[57]&P[56]&P[55]&P[54]&G[53]) | (P[57]&P[56]&P[55]&P[54]&P[53]&G[52]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&G[51]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&G[50]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&G[49]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&G[48]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&G[47]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&G[46]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&G[45]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&G[44]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&G[43]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[59] = G[58] | (P[58]&G[57]) | (P[58]&P[57]&G[56]) | (P[58]&P[57]&P[56]&G[55]) | (P[58]&P[57]&P[56]&P[55]&G[54]) | (P[58]&P[57]&P[56]&P[55]&P[54]&G[53]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&G[52]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&G[51]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&G[50]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&G[49]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&G[48]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&G[47]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&G[46]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&G[45]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&G[44]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&G[43]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[60] = G[59] | (P[59]&G[58]) | (P[59]&P[58]&G[57]) | (P[59]&P[58]&P[57]&G[56]) | (P[59]&P[58]&P[57]&P[56]&G[55]) | (P[59]&P[58]&P[57]&P[56]&P[55]&G[54]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&G[53]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&G[52]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&G[51]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&G[50]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&G[49]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&G[48]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&G[47]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&G[46]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&G[45]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&G[44]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&G[43]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[61] = G[60] | (P[60]&G[59]) | (P[60]&P[59]&G[58]) | (P[60]&P[59]&P[58]&G[57]) | (P[60]&P[59]&P[58]&P[57]&G[56]) | (P[60]&P[59]&P[58]&P[57]&P[56]&G[55]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&G[54]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&G[53]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&G[52]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&G[51]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&G[50]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&G[49]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&G[48]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&G[47]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&G[46]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&G[45]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&G[44]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&G[43]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[62] = G[61] | (P[61]&G[60]) | (P[61]&P[60]&G[59]) | (P[61]&P[60]&P[59]&G[58]) | (P[61]&P[60]&P[59]&P[58]&G[57]) | (P[61]&P[60]&P[59]&P[58]&P[57]&G[56]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&G[55]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&G[54]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&G[53]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&G[52]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&G[51]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&G[50]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&G[49]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&G[48]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&G[47]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&G[46]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&G[45]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&G[44]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&G[43]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign c[63] = G[62] | (P[62]&G[61]) | (P[62]&P[61]&G[60]) | (P[62]&P[61]&P[60]&G[59]) | (P[62]&P[61]&P[60]&P[59]&G[58]) | (P[62]&P[61]&P[60]&P[59]&P[58]&G[57]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&G[56]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&G[55]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&G[54]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&G[53]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&G[52]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&G[51]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&G[50]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&G[49]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&G[48]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&G[47]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&G[46]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&G[45]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&G[44]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&G[43]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);
assign Cout = G[63] | (P[63]&G[62]) | (P[63]&P[62]&G[61]) | (P[63]&P[62]&P[61]&G[60]) | (P[63]&P[62]&P[61]&P[60]&G[59]) | (P[63]&P[62]&P[61]&P[60]&P[59]&G[58]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&G[57]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&G[56]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&G[55]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&G[54]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&G[53]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&G[52]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&G[51]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&G[50]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&G[49]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&G[48]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&G[47]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&G[46]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&G[45]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&G[44]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&G[43]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&G[42]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&G[41]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&G[40]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&G[39]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&G[38]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&G[37]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&G[36]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&G[35]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&G[34]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&G[33]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&G[32]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&G[31]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&G[30]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&G[29]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&G[28]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&G[27]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[63]&P[62]&P[61]&P[60]&P[59]&P[58]&P[57]&P[56]&P[55]&P[54]&P[53]&P[52]&P[51]&P[50]&P[49]&P[48]&P[47]&P[46]&P[45]&P[44]&P[43]&P[42]&P[41]&P[40]&P[39]&P[38]&P[37]&P[36]&P[35]&P[34]&P[33]&P[32]&P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&c[0]);

endmodule